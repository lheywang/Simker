* Mixed-signal simulation: clk_div + counter
.control
  pre_osdi ./driver.osdi
.endc

* --- 1. BRIDGE MODELS ---
.model a2d adc_bridge(in_low=0.4 in_high=0.8)
.model d2a dac_bridge(out_low=0.0 out_high=1.0)

* --- 2. ANALOG SOURCES ---
Vclk clk_a 0 PULSE(0 1 0 1n 1n 100n 200n)
Vrst rst_a 0 PWL(0 0 450n 0 451n 1)

* --- 3. INPUT BRIDGES (Analog to Digital) ---
abridge_in [clk_a rst_a] [clk_d rst_d] a2d

* --- 4. DIGITAL COSIM INSTANCE ---
Atop [rst_d clk_d] [q3_d q2_d q1_d q0_d] top
.model top d_cosim simulation="./top.so"

* --- 5. OUTPUT BRIDGES (Digital to Analog) ---
abridge_out0 [q0_d] [q0_a] d2a
abridge_out1 [q1_d] [q1_a] d2a
abridge_out2 [q2_d] [q2_a] d2a
abridge_out3 [q3_d] [q3_a] d2a

* --- 6. ANALOG DRIVERS & LOADS ---
.Model driver_model driver
.subckt driver in out
  Ndriver in out driver_model
.ends

Xdrv0 q0_a o0 driver
Xdrv1 q1_a o1 driver
Xdrv2 q2_a o2 driver
Xdrv3 q3_a o3 driver

Rload0 o0 o0c 100
Rload1 o1 o1c 100
Rload2 o2 o2c 100
Rload3 o3 o3c 100

Cload0 o0c 0 1n
Cload1 o1c 0 1n
Cload2 o2c 0 1n
Cload3 o3c 0 1n

* --- 7. SIMULATION ---
.tran 10n 15u

.control
  run
  * Plot the analog clock and the final driver outputs
  plot v(clk_a) v(o3c)+24 v(o2c)+18 v(o1c)+12 v(o0c)+6 v(rst_a)-6
.endc
.end
